library IEEE;
use IEEE.std_logic_1164.all;

entity LUT is
port (
    F	:	in std_logic_vector(5 downto 0);
    A	: 	out std_logic_vector(35 downto 0)
    );
  end LUT;
  
  architecture tabla of LUT is
 begin
  process(F)
  begin case F is
	--when "000000" => A <= "000001100110011001100110011001100110"; 
	--when "000001" => A <= "111100110011001100110011001100110100"; 
	--when "000010" => A <= "010011001100110011001100110011001100"; 
	--when "000011" => A <= "111100110011001100110011001100110100"; 
	--when "000100" => A <= "000001100110011001100110011001100110";
	when "000000" => A <= "010000000000000000000000000000000000"; 
	when "000001" => A <= "010000000000000000000000000000000000"; 
	when "000010" => A <= "010000000000000000000000000000000000"; 
	when "000011" => A <= "010000000000000000000000000000000000"; 
	when "000100" => A <= "010000000000000000000000000000000000";
	when others => A <= (others => '0'); 

       end case;
    end process;
  end tabla;
